/**
 * Demultiplexor:
 * {a, b} = {in, 0} if sel == 0
 *          {0, in} if sel == 1
 */

`default_nettype none
module DMux(
    input in,
    input sel,
    output a,
    output b
);

    // No need to implement this chip
    assign a = ~sel&in;
    assign b = sel&in;

endmodule
