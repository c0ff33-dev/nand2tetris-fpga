/**
 * 4-way demultiplexor:
 * {a, b, c, d} = {in, 0, 0, 0} if sel == 00
 *                {0, in, 0, 0} if sel == 01
 *                {0, 0, in, 0} if sel == 10
 *                {0, 0, 0, in} if sel == 11
 */

`default_nettype none
module DMux4Way(
	input in,
	input [1:0] sel,
    output a,
	output b,
	output c,
	output d
);
	
	// Put your code here:
	assign a = (sel==0) ? in : 0;
	assign b = (sel==1) ? in : 0;
	assign c = (sel==2) ? in : 0;
	assign d = (sel==3) ? in : 0;

endmodule