/**
 * 16 bit bitwise And:
 * for i = 0..15: out[i] = (a[i] and b[i])
 */

`default_nettype none
module And16(
    input [15:0] a,
    input [15:0] b,
    output [15:0] out
);

    // Put your code here:
    assign out = a&b; // bitwise AND (verilog primitive)

endmodule
