/**
 * Buffer:
 * out = in
 */

`default_nettype none
module Buffer(
	input in,
	output out
);

	assign out = in; // combinatorial memory

endmodule
