/**
 * Buffer:
 * out = in
 */

`default_nettype none
module Buffer(
	input in,
	output out
);

	// No need to implement this chip
	assign out = in;

endmodule
