/**
 * 16-bit bitwise Or:
 * for i = 0..15: out[i] = (a[i] or b[i])
 */

`default_nettype none
module Or16(
	input [15:0] a,
	input [15:0] b,
	output [15:0] out
);

	assign out = a|b; // bitwise OR

endmodule
