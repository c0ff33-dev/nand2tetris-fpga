 /**
 * Or gate:
 * out = 1 if (a == 1 or b == 1)
 *       0 otherwise
 */

`default_nettype none
module Or(
	input a,
	input b,
	output out
);

	// Put your code here:
	or(out,a,b); // bitwise OR (verilog primitive)

endmodule
