/**
 * Adds two 16 bit values.
 * The most significant carry bit is ignored.
 * out = a + b (16 bit)
 */

`default_nettype none
module Add16(
	input [15:0] a,
	input [15:0] b,
	output [15:0] out
);

	// Put your code here:
	assign out = a + b;

endmodule
