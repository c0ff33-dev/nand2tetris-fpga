/**
 * 1 bit register:
 * If load[t] == 1 then out[t+1] = in[t]
 *    else out does not change (out[t+1] = out[t])
 */

`default_nettype none
module Bit(
    input clk,
    input in,
    input load,
    output reg out = 0
);

    // No need to implement this chip
    always @(posedge clk)
        out <= load?in:out;

endmodule
